interface mux_intf ();
  logic din_0,din_1,din_2,din_3;
  logic y;
  logic[1:0] sel;  
  endinterface
