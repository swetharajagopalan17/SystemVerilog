interface intf_seq (input logic clock ,reset);
  logic in_d ;
  logic dout ;
  
endinterface
