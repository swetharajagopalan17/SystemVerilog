class transaction;
  rand bit j;
  rand bit k;
  //clk and reset are top level so no need to declare here 
  bit q;
  
  //define constraints here 
  
  //printing stuff 
  
  
endclass
