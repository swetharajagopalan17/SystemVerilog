class transaction ;
  rand bit Din ;
  bit dout ;
endclass
