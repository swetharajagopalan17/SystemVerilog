class config_db;
  static mailbox gen2driv_mb = new();
  static mailbox mon2sb_mb = new();
endclass
