interface jk_intf(input logic clk);
  logic j;
  logic k;
  logic q;
endinterface
