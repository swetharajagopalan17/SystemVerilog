class transaction ;
  
  rand bit j,k;
  bit qout;
 
endclass
