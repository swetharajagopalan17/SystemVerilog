interface jk_ff_intf (input logic clk);
  
  logic j,k;
  logic qout;
  
 endinterface
